module test_clint_detailed;
    reg clk;
    reg rst_n;
    reg bus_en;
    reg bus_we;
    reg [31:0] bus_addr;
    reg [31:0] bus_wdata;
    wire [31:0] bus_rdata;
    wire bus_ready;
    wire timer_irq;
    wire software_irq;
    
    // 实例化CLINT
    clint u_clint (
        .clk(clk),
        .rst_n(rst_n),
        .bus_en(bus_en),
        .bus_we(bus_we),
        .bus_addr(bus_addr),
        .bus_wdata(bus_wdata),
        .bus_rdata(bus_rdata),
        .bus_ready(bus_ready),
        .timer_irq_o(timer_irq),
        .software_irq_o(software_irq),
        .irq_enable(1'b1),
        .timer_mode(2'b00)  // 周期性模式
    );
    
    // 时钟生成
    always #5 clk = ~clk;
    
    // 测试任务：写入寄存器
    task write_reg;
        input [31:0] addr;
        input [31:0] data;
        begin
            @(posedge clk);
            bus_en = 1'b1;
            bus_we = 1'b1;
            bus_addr = addr;
            bus_wdata = data;
            @(posedge clk);
            while (!bus_ready) @(posedge clk);
            bus_en = 1'b0;
            bus_we = 1'b0;
            #10;
            $display("[%0t] 写入寄存器 0x%08h = 0x%08h", $time, addr, data);
        end
    endtask
    
    // 测试任务：读取寄存器
    task read_reg;
        input [31:0] addr;
        output [31:0] data;
        begin
            @(posedge clk);
            bus_en = 1'b1;
            bus_we = 1'b0;
            bus_addr = addr;
            @(posedge clk);
            while (!bus_ready) @(posedge clk);
            data = bus_rdata;
            bus_en = 1'b0;
            #10;
            $display("[%0t] 读取寄存器 0x%08h = 0x%08h", $time, addr, data);
        end
    endtask
    
    // 监控定时器值
    task monitor_timer;
        integer i;
        begin
            for (i = 0; i < 10; i = i + 1) begin
                #100;  // 每100个时间单位检查一次
                begin
                    reg [31:0] mtime_low, mtime_high, mtimecmp_low;
                    read_reg(32'h0200BFF8, mtime_low);
                    read_reg(32'h0200BFFC, mtime_high);
                    read_reg(32'h02004000, mtimecmp_low);
                    $display("[%0t] MTIME=0x%08h_%08h, MTIMECMP低32位=0x%08h, timer_irq=%b", 
                             $time, mtime_high, mtime_low, mtimecmp_low, timer_irq);
                end
            end
        end
    endtask
    
    initial begin
        $dumpfile("clint_detailed_test.vcd");
        $dumpvars(0, test_clint_detailed);
        
        // 初始化
        clk = 0;
        rst_n = 0;
        bus_en = 0;
        bus_we = 0;
        bus_addr = 0;
        bus_wdata = 0;
        
        // 复位
        #20 rst_n = 1;
        
        $display("=== CLINT 详细测试开始 ===");
        $display("时钟频率: 100MHz (周期10ns)");
        
        // 测试1：检查定时器是否在运行
        $display("\n测试1：检查定时器基础功能");
        begin
            reg [31:0] mtime1, mtime2;
            read_reg(32'h0200BFF8, mtime1);
            #100;  // 等待10个时钟周期
            read_reg(32'h0200BFF8, mtime2);
            if (mtime2 > mtime1) 
                $display("  ✅ 定时器正在运行: %d -> %d", mtime1, mtime2);
            else
                $display("  ❌ 定时器没有运行: %d -> %d", mtime1, mtime2);
        end
        
        // 测试2：定时器中断
        $display("\n测试2：定时器中断测试");
        
        // 读取当前定时器值
        begin
            reg [31:0] current_mtime;
            read_reg(32'h0200BFF8, current_mtime);
            $display("  当前MTIME低32位: 0x%08h (%0d)", current_mtime, current_mtime);
        end
        
        // 设置定时器比较值为当前值+10
        begin
            reg [31:0] current_mtime;
            read_reg(32'h0200BFF8, current_mtime);
            write_reg(32'h02004000, current_mtime + 10);
            $display("  设置MTIMECMP = 当前值 + 10");
        end
        
        // 监控一段时间
        $display("\n  监控定时器10个周期...");
        monitor_timer();
        
        // 检查中断是否触发
        if (timer_irq) begin
            $display("  ✅ 定时器中断成功触发");
            
            // 测试周期性模式：清除中断后应该再次触发
            $display("\n  测试周期性模式...");
            #200;
            
            if (timer_irq) 
                $display("  ✅ 周期性中断工作正常");
            else
                $display("  ⚠️  周期性中断可能有问题");
                
        end else begin
            $display("  ❌ 定时器中断没有触发");
            
            // 诊断：检查寄存器值
            begin
                reg [31:0] mtime_low, mtime_high, mtimecmp_low, mtimecmp_high;
                read_reg(32'h0200BFF8, mtime_low);
                read_reg(32'h0200BFFC, mtime_high);
                read_reg(32'h02004000, mtimecmp_low);
                read_reg(32'h02004004, mtimecmp_high);
                
                $display("  诊断信息:");
                $display("    MTIME: 0x%08h_%08h (%0d)", mtime_high, mtime_low, {mtime_high, mtime_low});
                $display("    MTIMECMP: 0x%08h_%08h (%0d)", mtimecmp_high, mtimecmp_low, {mtimecmp_high, mtimecmp_low});
                $display("    差值: %0d", ({mtime_high, mtime_low} - {mtimecmp_high, mtimecmp_low}));
                $display("    中断使能: 1 (固定)");
            end
        end
        
        // 测试3：软件中断
        $display("\n测试3：软件中断测试");
        write_reg(32'h02000000, 32'h1);  // 触发软件中断
        #10;
        if (software_irq) $display("  ✅ 软件中断触发成功");
        else $display("  ❌ 软件中断失败");
        
        write_reg(32'h02000000, 32'h0);  // 清除软件中断
        #10;
        if (!software_irq) $display("  ✅ 软件中断清除成功");
        else $display("  ❌ 软件中断清除失败");
        
        $display("\n=== CLINT 详细测试完成 ===");
        
        #100 $finish;
    end
    
    // 监视中断信号
    always @(posedge timer_irq) begin
        $display("[%0t] ⏰ 定时器中断触发!", $time);
    end
    
    always @(posedge software_irq) begin
        $display("[%0t] 🖥️  软件中断触发!", $time);
    end
    
endmodule